// mem controller init file
